//--------------------------------------------------------------------
// Author: Lalit Prasad Peri (lalitprasad@vt.edu)
// Group5 Project: Advance VLSI Design, ECE5545 Spring2024 
//--------------------------------------------------------------------
// Simple Verilog TB for Synthesis
//--------------------------------------------------------------------

module testbench(

 input aclk,
 input aresetn,
 input srst,

 input mst0_aclk,
 input mst1_aclk,
 input mst2_aclk,
 input mst3_aclk,

 input slv0_aclk,
 input slv1_aclk,
 input slv2_aclk,
 input slv3_aclk,

 input  slv0_awvalid,
 input  slv0_wvalid,
 input  slv0_arvalid,
 input  slv1_awvalid,
 input  slv1_wvalid,
 input  slv1_arvalid,
 input  slv2_awvalid,
 input  slv2_wvalid,
 input  slv2_arvalid,
 input  slv3_awvalid,
 input  slv3_wvalid,
 input  slv3_arvalid,
 input  mst0_bvalid,
 input  mst0_rvalid,
 input  mst1_bvalid,
 input  mst1_rvalid,
 input  mst2_bvalid,
 input  mst2_rvalid,
 input  mst3_bvalid,
 input  mst3_rvalid,
 input  slv0_bready,
 input  slv0_rready,
 input  slv1_bready,
 input  slv1_rready,
 input  slv2_bready,
 input  slv2_rready,
 input  slv3_bready,
 input  slv3_rready,
 input  mst0_awready,
 input  mst0_wready,
 input  mst0_arready,
 input  mst1_awready,
 input  mst1_wready,
 input  mst1_arready,
 input  mst2_awready,
 input  mst2_wready,
 input  mst2_arready,
 input  mst3_awready,
 input  mst3_wready,
 input  mst3_arready,
 output slv0_bvalid,
 output slv0_rvalid,
 output slv1_bvalid,
 output slv1_rvalid,
 output slv2_bvalid,
 output slv2_rvalid,
 output slv3_bvalid,
 output slv3_rvalid,
 output mst0_awvalid,
 output mst0_wvalid,
 output mst0_arvalid,
 output mst1_awvalid,
 output mst1_wvalid,
 output mst1_arvalid,
 output mst2_awvalid,
 output mst2_wvalid,
 output mst2_arvalid,
 output mst3_awvalid,
 output mst3_wvalid,
 output mst3_arvalid,
 output slv0_awready,
 output slv0_wready,
 output slv0_arready,
 output slv1_awready,
 output slv1_wready,
 output slv1_arready,
 output slv2_awready,
 output slv2_wready,
 output slv2_arready,
 output slv3_awready,
 output slv3_wready,
 output slv3_arready,
 output mst0_bready,
 output mst0_rready,
 output mst1_bready,
 output mst1_rready,
 output mst2_bready,
 output mst2_rready,
 output mst3_bready,
 output mst3_rready 

);

//DUT
axicb_crossbar_top axicb_crossbar_top (

        .aclk         (aclk),    
        .aresetn      (aresetn),
        .srst         (srst),    

        .mst0_aclk      (mst0_aclk),
        .mst0_aresetn   (aresetn), 
        .mst0_srst      (srst),     
        .mst1_aclk      (mst1_aclk),
        .mst1_aresetn   (aresetn), 
        .mst1_srst      (srst),     
        .mst2_aclk      (mst2_aclk),
        .mst2_aresetn   (aresetn), 
        .mst2_srst      (srst),     
        .mst3_aclk      (mst3_aclk),
        .mst3_aresetn   (aresetn), 
        .mst3_srst      (srst),     

        .slv0_aclk      (slv0_aclk),
        .slv0_aresetn   (aresetn), 
        .slv0_srst      (srst),     
        .slv1_aclk      (slv1_aclk),
        .slv1_aresetn   (aresetn), 
        .slv1_srst      (srst),     
        .slv2_aclk      (slv2_aclk),
        .slv2_aresetn   (aresetn), 
        .slv2_srst      (srst),     
        .slv3_aclk      (slv3_aclk),
        .slv3_aresetn   (aresetn), 
        .slv3_srst      (srst),     

        .slv0_awvalid   (slv0_awvalid), 
        .slv0_wvalid    (slv0_wvalid), 
        .slv0_arvalid   (slv0_arvalid), 
        .slv1_awvalid   (slv1_awvalid), 
        .slv1_wvalid    (slv1_wvalid), 
        .slv1_arvalid   (slv1_arvalid), 
        .slv2_awvalid   (slv2_awvalid), 
        .slv2_wvalid    (slv2_wvalid), 
        .slv2_arvalid   (slv2_arvalid), 
        .slv3_awvalid   (slv3_awvalid), 
        .slv3_wvalid    (slv3_wvalid), 
        .slv3_arvalid   (slv3_arvalid), 
        .mst0_bvalid    (mst0_bvalid), 
        .mst0_rvalid    (mst0_rvalid), 
        .mst1_bvalid    (mst1_bvalid), 
        .mst1_rvalid    (mst1_rvalid), 
        .mst2_bvalid    (mst2_bvalid), 
        .mst2_rvalid    (mst2_rvalid), 
        .mst3_bvalid    (mst3_bvalid), 
        .mst3_rvalid    (mst3_rvalid), 
        .slv0_bready    (slv0_bready), 
        .slv0_rready    (slv0_rready), 
        .slv1_bready    (slv1_bready), 
        .slv1_rready    (slv1_rready), 
        .slv2_bready    (slv2_bready), 
        .slv2_rready    (slv2_rready), 
        .slv3_bready    (slv3_bready), 
        .slv3_rready    (slv3_rready), 
        .mst0_awready   (mst0_awready), 
        .mst0_wready    (mst0_wready), 
        .mst0_arready   (mst0_arready), 
        .mst1_awready   (mst1_awready), 
        .mst1_wready    (mst1_wready), 
        .mst1_arready   (mst1_arready), 
        .mst2_awready   (mst2_awready), 
        .mst2_wready    (mst2_wready), 
        .mst2_arready   (mst2_arready), 
        .mst3_awready   (mst3_awready), 
        .mst3_wready    (mst3_wready), 
        .mst3_arready   (mst3_arready), 
        .slv0_bvalid    (slv0_bvalid), 
        .slv0_rvalid    (slv0_rvalid), 
        .slv1_bvalid    (slv1_bvalid), 
        .slv1_rvalid    (slv1_rvalid), 
        .slv2_bvalid    (slv2_bvalid), 
        .slv2_rvalid    (slv2_rvalid), 
        .slv3_bvalid    (slv3_bvalid), 
        .slv3_rvalid    (slv3_rvalid), 
        .mst0_awvalid   (mst0_awvalid), 
        .mst0_wvalid    (mst0_wvalid), 
        .mst0_arvalid   (mst0_arvalid), 
        .mst1_awvalid   (mst1_awvalid), 
        .mst1_wvalid    (mst1_wvalid), 
        .mst1_arvalid   (mst1_arvalid), 
        .mst2_awvalid   (mst2_awvalid), 
        .mst2_wvalid    (mst2_wvalid), 
        .mst2_arvalid   (mst2_arvalid), 
        .mst3_awvalid   (mst3_awvalid), 
        .mst3_wvalid    (mst3_wvalid), 
        .mst3_arvalid   (mst3_arvalid), 
        .slv0_awready   (slv0_awready), 
        .slv0_wready    (slv0_wready), 
        .slv0_arready   (slv0_arready), 
        .slv1_awready   (slv1_awready), 
        .slv1_wready    (slv1_wready), 
        .slv1_arready   (slv1_arready), 
        .slv2_awready   (slv2_awready), 
        .slv2_wready    (slv2_wready), 
        .slv2_arready   (slv2_arready), 
        .slv3_awready   (slv3_awready), 
        .slv3_wready    (slv3_wready), 
        .slv3_arready   (slv3_arready), 
        .mst0_bready    (mst0_bready), 
        .mst0_rready    (mst0_rready), 
        .mst1_bready    (mst1_bready), 
        .mst1_rready    (mst1_rready), 
        .mst2_bready    (mst2_bready), 
        .mst2_rready    (mst2_rready), 
        .mst3_bready    (mst3_bready), 
        .mst3_rready    (mst3_rready),  

        // Master Agent 0 interface
        .slv0_awaddr  ('h0),
        .slv0_awprot  ('h0),
        .slv0_awid    ('h0),
        .slv0_awuser  ('h0),
        .slv0_wdata   ('h0),
        .slv0_wstrb   ('h0),
        .slv0_wuser   ('h0),
        .slv0_araddr  ('h0),
        .slv0_arprot  ('h0),
        .slv0_arid    ('h0),
        .slv0_aruser  ('h0),
        .slv0_bid     (), 
        .slv0_bresp   (),
        .slv0_buser   (),
        .slv0_rid     (),
        .slv0_rresp   (),
        .slv0_rdata   (),
        .slv0_ruser   (),
        // Master Agent 1 interface
        .slv1_awaddr  ('h0),
        .slv1_awprot  ('h0),
        .slv1_awid    ('h0),
        .slv1_awuser  ('h0),
        .slv1_wdata   ('h0),
        .slv1_wstrb   ('h0),
        .slv1_wuser   ('h0),
        .slv1_araddr  ('h0),
        .slv1_arprot  ('h0),
        .slv1_arid    ('h0),
        .slv1_aruser  ('h0),
        .slv1_bid     (), 
        .slv1_bresp   (),
        .slv1_buser   (),
        .slv1_rid     (),
        .slv1_rresp   (),
        .slv1_rdata   (),
        .slv1_ruser   (),
        // Master Agent 2 interface
        .slv2_awaddr  ('h0),
        .slv2_awprot  ('h0),
        .slv2_awid    ('h0),
        .slv2_awuser  ('h0),
        .slv2_wdata   ('h0),
        .slv2_wstrb   ('h0),
        .slv2_wuser   ('h0),
        .slv2_araddr  ('h0),
        .slv2_arprot  ('h0),
        .slv2_arid    ('h0),
        .slv2_aruser  ('h0),
        .slv2_bid     (), 
        .slv2_bresp   (),
        .slv2_buser   (),
        .slv2_rid     (),
        .slv2_rresp   (),
        .slv2_rdata   (),
        .slv2_ruser   (),
        // Master Agent 3 interface
        .slv3_awaddr  ('h0),
        .slv3_awprot  ('h0),
        .slv3_awid    ('h0),
        .slv3_awuser  ('h0),
        .slv3_wdata   ('h0),
        .slv3_wstrb   ('h0),
        .slv3_wuser   ('h0),
        .slv3_araddr  ('h0),
        .slv3_arprot  ('h0),
        .slv3_arid    ('h0),
        .slv3_aruser  ('h0),
        .slv3_bid     (), 
        .slv3_bresp   (),
        .slv3_buser   (),
        .slv3_rid     (),
        .slv3_rresp   (),
        .slv3_rdata   (),
        .slv3_ruser   (),

        // Slave Agent 0 interface
        .mst0_bid     ('h0),
        .mst0_bresp   ('h0),
        .mst0_buser   ('h0),
        .mst0_rid     ('h0),
        .mst0_rresp   ('h0),
        .mst0_rdata   ('h0),
        .mst0_ruser   ('h0),
        .mst0_awaddr  (),
        .mst0_awprot  (),
        .mst0_awid    (),
        .mst0_awuser  (),
        .mst0_wdata   (),
        .mst0_wstrb   (),
        .mst0_wuser   (),
        .mst0_araddr  (),
        .mst0_arprot  (),
        .mst0_arid    (),
        .mst0_aruser  (),
        // Slave Agent 1 interface
        .mst1_bid     ('h0),
        .mst1_bresp   ('h0),
        .mst1_buser   ('h0),
        .mst1_rid     ('h0),
        .mst1_rresp   ('h0),
        .mst1_rdata   ('h0),
        .mst1_ruser   ('h0),
        .mst1_awaddr  (),
        .mst1_awprot  (),
        .mst1_awid    (),
        .mst1_awuser  (),
        .mst1_wdata   (),
        .mst1_wstrb   (),
        .mst1_wuser   (),
        .mst1_araddr  (),
        .mst1_arprot  (),
        .mst1_arid    (),
        .mst1_aruser  (),
        // Slave Agent 2 interface
        .mst2_bid     ('h0),
        .mst2_bresp   ('h0),
        .mst2_buser   ('h0),
        .mst2_rid     ('h0),
        .mst2_rresp   ('h0),
        .mst2_rdata   ('h0),
        .mst2_ruser   ('h0),
        .mst2_awaddr  (),
        .mst2_awprot  (),
        .mst2_awid    (),
        .mst2_awuser  (),
        .mst2_wdata   (),
        .mst2_wstrb   (),
        .mst2_wuser   (),
        .mst2_araddr  (),
        .mst2_arprot  (),
        .mst2_arid    (),
        .mst2_aruser  (),
        // Slave Agent 3 interface
        .mst3_bid     ('h0),
        .mst3_bresp   ('h0),
        .mst3_buser   ('h0),
        .mst3_rid     ('h0),
        .mst3_rresp   ('h0),
        .mst3_rdata   ('h0),
        .mst3_ruser   ('h0),
        .mst3_awaddr  (),
        .mst3_awprot  (),
        .mst3_awid    (),
        .mst3_awuser  (),
        .mst3_wdata   (),
        .mst3_wstrb   (),
        .mst3_wuser   (),
        .mst3_araddr  (),
        .mst3_arprot  (),
        .mst3_arid    (),
        .mst3_aruser  () 

    );

//--------------------------------------------------------------------
endmodule


